`timescale 1ns / 1ps


module hexto7segment(
    input [15:0] x,
    output reg [7:0] r1,
    output reg [7:0] r2,
    output reg [7:0] r3,
    output reg [7:0] r4
    );
    
    always @(*)begin
        case(x/1000)
            16'h0: r4 = 8'b00000011;
            16'h1 : r4 = 8'b10011111;
            16'h2 : r4 = 8'b00100101;
            16'h3 : r4 = 8'b00001101;
            16'h4 : r4 = 8'b10011001;
            16'h5 : r4 = 8'b01001001;
            16'h6 : r4 = 8'b01000001;
            16'h7 : r4 = 8'b00011111;
            16'h8 : r4 = 8'b00000001;
            16'h9 : r4 = 8'b00011001;
       endcase
       case((x/100)%10)
            16'h0: r3 = 8'b00000010;
            16'h1 : r3 = 8'b10011110;
            16'h2 : r3 = 8'b00100100;
            16'h3 : r3 = 8'b00001100;
            16'h4 : r3 = 8'b10011000;
            16'h5 : r3 = 8'b01001000;
            16'h6 : r3 = 8'b01000000;
            16'h7 : r3 = 8'b00011110;
            16'h8 : r3 = 8'b00000000;
            16'h9 : r3 = 8'b00011000;
       endcase
       case((x/10)%10)
            16'h0: r2 = 8'b00000011;
            16'h1 : r2 = 8'b10011111;
            16'h2 : r2 = 8'b00100101;
            16'h3 : r2 = 8'b00001101;
            16'h4 : r2 = 8'b10011001;
            16'h5 : r2 = 8'b01001001;
            16'h6 : r2 = 8'b01000001;
            16'h7 : r2 = 8'b00011111;
            16'h8 : r2 = 8'b00000001;
            16'h9 : r2 = 8'b00011001;
       endcase
       case(x%10)
            16'd0: r1 = 8'b00000011;
            16'd1 : r1 = 8'b10011111;
            16'd2 : r1 = 8'b00100101;
            16'd3 : r1 = 8'b00001101;
            16'd4 : r1 = 8'b10011001;
            16'd5 : r1 = 8'b01001001;
            16'd6 : r1 = 8'b01000001;
            16'd7 : r1 = 8'b00011111;
            16'd8 : r1 = 8'b00000001;
            16'd9 : r1 = 8'b00011001;
       endcase
       end
endmodule
